`timescale 1ns / 1p
module FA_FSM(
		input clk,
		input reset,
		input wd_selec,
		input write_en,
		input [1:0] read_add1,
		input [1:0] read_add2,
		input [1:0] write_add,
		output is_zero,
		output [31:0] result
    );

	

endmodule
